module decoder ( input wire [4:0] x, output reg [6:0] y );

    always @(x) begin
        case(x)
            'd0:     y <= 'b1000000;        // 0, O
            'd1:     y <= 'b1111001;        // 1
            'd2:     y <= 'b0100100;        // 2
            'd3:     y <= 'b0110000;        // 3
            'd4:     y <= 'b0011001;        // 4
            'd5:     y <= 'b0010010;        // 5, S
            'd6:     y <= 'b0000010;        // 6
            'd7:     y <= 'b1111000;        // 7
            'd8:     y <= 'b0000000;        // 8
            'd9:     y <= 'b0010000;        // 9
            'd10:    y <= 'b0001000;        // A
            'd11:    y <= 'b0000011;        // B
            'd12:    y <= 'b1000110;        // C
            'd13:    y <= 'b0100001;        // D
            'd14:    y <= 'b0000110;        // E
            'd15:    y <= 'b0001110;        // F
            'd16:    y <= 'b0101111;        // r
            default: y <= 'b1111111;
        endcase
    end

endmodule